----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/18/2022 12:56:11 PM
-- Design Name: 
-- Module Name: player - player_1
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity player is
   Port ( 
      clk, reset: in std_logic;
      btn: in std_logic_vector(3 downto 0);
      video_on: in std_logic;
      pixel_x, pixel_y: in std_logic_vector(9 downto 0);
      graph_rgb: out std_logic_vector(2 downto 0);
      doing_assignment: out std_logic;
      holding_breath: out std_logic;
      blocking_view: out std_logic;
      blocking_door: out std_logic
   );
end player;

architecture player_1 of player is
   type player_face is array(0 to 30) of std_logic_vector(0 to 30); -- Face is 31x31 pixels.
   constant HAPPY_ROM: player_face := (
      "0000000000001111111000000000000",
      "0000000001110000000111000000000",
      "0000000110000000000000110000000",
      "0000001000000000000000001000000",
      "0000010000000000000000000100000",
      "0000100000000000000000000010000",
      "0001000000000000000000000001000",
      "0010000001110000001110000000100",
      "0010000001110000001110000000100",
      "0100000001110000001110000000010",
      "0100000000000000000000000000010",
      "0100000000000000000000000000010",
      "1000000000000000000000000000001",
      "1000000000000000000000000000001",
      "1000000000000000000000000000001",
      "1000000000000000000000000000001",
      "1000000000000000000000000000001",
      "1000000000000000000000000000001",
      "1000000000000000000000000000001",
      "0100000001000000000001000000010",
      "0100000000100000000010000000010",
      "0100000000010000000100000000010",
      "0010000000001000001000000000100",
      "0010000000000111110000000000100",
      "0001000000000000000000000001000",
      "0000100000000000000000000010000",
      "0000010000000000000000000100000",
      "0000001000000000000000001000000",
      "0000000110000000000000110000000",
      "0000000001110000000111000000000",
      "0000000000001111111000000000000"
      );
   constant LOSE_ROM: player_face := (
      "0000000000001111111000000000000",
      "0000000001110000000111000000000",
      "0000000110000000000000110000000",
      "0000001000000000000000001000000",
      "0000010000000000000000000100000",
      "0000100000000000000000000010000",
      "0001000000000000000000000001000",
      "0010000001110000001110000000100",
      "0010000001110000001110000000100",
      "0100000001110000001110000000010",
      "0100000000000000000000000000010",
      "0100000000000000000000000000010",
      "1000000000000000000000000000001",
      "1000000000000000000000000000001",
      "1000000000000000000000000000001",
      "1000000000000011100000000000001",
      "1000000000000100010000000000001",
      "1000000000001000001000000000001",
      "1000000000010000000100000000001",
      "0100000000010000000100000000010",
      "0100000000010000000100000000010",
      "0100000000010000000100000000010",
      "0010000000001000001000000000100",
      "0010000000000100010000000000100",
      "0001000000000011100000000001000",
      "0000100000000000000000000010000",
      "0000010000000000000000000100000",
      "0000001000000000000000001000000",
      "0000000110000000000000110000000",
      "0000000001110000000111000000000",
      "0000000000001111111000000000000"
      );
   constant SCARED_ROM: player_face := (
      "0000000000001111111000000000000",
      "0000000001110000000111000000000",
      "0000000110000000000000110000000",
      "0000001000000000000000001000000",
      "0000010000000000000000000100000",
      "0000100000000000000000000010000",
      "0001000000000000000000000001000",
      "0010000001110000001110000000100",
      "0010000001110000001110000000100",
      "0100000001110000001110000000010",
      "0100000010000000000000000000010",
      "0100000110000000000000000000010",
      "1000000110000000000000000000001",
      "1000000110000000000000000000001",
      "1000000110000000000000000000001",
      "1000000110000000000000000000001",
      "1000000100000000000000000000001",
      "1000000000000000000000000000001",
      "1000000000000000000000000000001",
      "0100000000000000000000000000010",
      "0100000000000000000000000000010",
      "0100000000000000000000000000010",
      "0010000000111111111100000000100",
      "0010000000000000000000000000100",
      "0001000000000000000000000001000",
      "0000100000000000000000000010000",
      "0000010000000000000000000100000",
      "0000001000000000000000001000000",
      "0000000110000000000000110000000",
      "0000000001110000000111000000000",
      "0000000000001111111000000000000"
      );
   type assignment is array(0 to 12) of std_logic_vector(0 to 14); --paper & pencil is 13x15
   constant assignment_ROM: assignment := (
      "000001111111111",
      "000001000000001",
      "000001000000001",
      "000011011101101",
      "000101000000001",
      "001001010110101",
      "010001000000001",
      "100001011100001",
      "000001000000001",
      "000001000000001",
      "000001000000001",
      "000001000000001",
      "000001111111111"
      );
   type hand is array(0 to 19) of std_logic_vector(0 to 9); --hand is 20x10
   constant hand_ROM: hand := (
      "0000010000",
      "0011010000",
      "0001010100",
      "0001010101",
      "1001111101",
      "1011000110",
      "0110000010",
      "0010000010",
      "0010000010",
      "0010000010",
      "0010000010",
      "0001000100",
      "0001000100",
      "0001000100",
      "0001000100",
      "0001000100",
      "0001000100",
      "0001000100",
      "0001000100",
      "0001000100"
   );
   
   type backpack is array(0 to 15) of std_logic_vector(0 to 8); --backpack is 16x9
   constant backpack_ROM: backpack := (
      "111100000",
      "111111000",
      "110111100",
      "110011100",
      "100001110",
      "100000111",
      "101000011",
      "101000011",
      "101000011",
      "101000011",
      "100000011",
      "100000011",
      "110000111",
      "110000111",
      "111111110",
      "111111100"
   );
begin


end player_1;
